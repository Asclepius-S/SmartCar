`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:48:26 06/26/2019 
// Design Name: 
// Module Name:    SEG7_LUT 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SEG7_LUT(dig,seg);
//////////////////////////////////////////////////////////////////////////////////
//		# 	DIG		seg 	    ____a____
//		1	1 OR I	1111001	 |		   |
//		2	2     	0100100	 f		   b
//		3	3		   0110000	 |		   |
//		4	4		   0011001	 ____g____
//		5	5 OR S	0010010	 |			|
//		6	6			0000010	 e		   c
//		7	7			1111000	 |		   |
//		8	8			0000000	 ____d____
//		9	9			0011000
//		0	0			1000000
//		10	p			0001000
//		11	a 			0001000
//		12	u OR w	1000001
//		13	e 			0000110
//		14	r			1001110
//		15	close		1111111
//////////////////////////////////////////////////////////////////////////////////
	input [3:0] dig;
	output reg [6:0] seg;

	always @ (dig)
	begin
		case(dig)
		4'h1: seg = 7'b1111001;//i
		4'h2: seg = 7'b0100100;
		4'h3: seg = 7'b0110000;
		4'h4: seg = 7'b0011001;
		4'h5: seg = 7'b0010010;//s
		4'h6: seg = 7'b0000010;
		4'h7: seg = 7'b1111000;
		4'h8: seg = 7'b0000000;
		4'h9: seg = 7'b0011000;
		4'h0: seg = 7'b1000000;
		4'ha: seg = 7'b0001000;//A
		4'hb: seg = 7'b0000011;//P
		4'hc: seg = 7'b1000110;//M
		4'hd: seg = 7'b0100001;//L
		4'he: seg = 7'b0000100;//F
		4'hf: seg = 7'b1111111;//close
		endcase
	end

endmodule

